----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/14/2023 10:54:55 PM
-- Design Name: 
-- Module Name: RCA_4 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ADD_SUB is
    Port ( A0 : in STD_LOGIC;
           A1 : in STD_LOGIC;
           A2 : in STD_LOGIC;
           A3 : in STD_LOGIC;
           M  : in STD_LOGIC;
           B0 : in STD_LOGIC;
           B1 : in STD_LOGIC;
           B2 : in STD_LOGIC;
           B3 : in STD_LOGIC;
           --C_in : in STD_LOGIC;
           S0 : out STD_LOGIC;
           S1 : out STD_LOGIC;
           S2 : out STD_LOGIC;
           S3 : out STD_LOGIC;
           --C_out : out STD_LOGIC;
           V : out STD_LOGIC;   --Overflow
           Zero : out STD_LOGIC );
end ADD_SUB;

architecture Behavioral of ADD_SUB is
component FA
     port (
     A: in std_logic;
     B: in std_logic;
     C_in: in std_logic;
     S: out std_logic;
     C_out: out std_logic);
 end component;

SIGNAL FA0_C, FA1_C, FA2_C, FA3_C, FA0_S, FA1_S, FA2_S, FA3_S  : std_logic;
SIGNAL B0_temp, B1_temp, B2_temp, B3_temp  : std_logic;
SIGNAL C_temp : std_logic;

begin
 FA_0 : FA
    port map (
    A => A0,
    B => B0_temp,
    C_in => M, 
    S => FA0_S,
    C_Out => FA0_C);   
 FA_1 : FA
    port map (
    A => A1,
    B => B1_temp,
    C_in => FA0_C,
    S => FA1_S,
    C_Out => FA1_C);
 FA_2 : FA
    port map (
    A => A2,
    B => B2_temp,
    C_in => FA1_C,
    S => FA2_S,
    C_Out => FA2_C);
 FA_3 : FA
    port map (
    A => A3,
    B => B3_temp,
    C_in => FA2_C,
    S => FA3_S,
    C_Out => C_temp);
         
B0_temp <= B0 XOR M;
B1_temp <= B1 XOR M;
B2_temp <= B2 XOR M;
B3_temp <= B3 XOR M;

S0 <= FA0_S;
S1 <= FA1_S;
S2 <= FA2_S;
S3 <= FA3_S;

V <= C_temp XOR FA2_C;
--C_out <= C_temp;
Zero <= NOT (FA0_S OR FA1_S OR FA2_S OR FA3_S);
  
end Behavioral;
